*                1 - Input A 2 - Input B 3 - VDD 5 - Output  
.subckt nor_gate 1 2 3 5 
.param ln = 1u wn = 1u

xmp1 4 1 3 3 pmos1v l=ln w= wn
xmp2 5 2 4 4 pmos1v l=ln w= wn

xmn1 5 1 0 0 nmos1v l=ln w= wn
xmn2 5 2 0 0 nmos1v l=ln w= wn
.ends
