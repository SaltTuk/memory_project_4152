[aimspice]
[description]
233
Ex3b
.include C:\Users\itsom\Desktop\FALL2022\TFE4152\90_nm_gpdk\gpdk90nm_ff.cir
.plot id(m:mn2:1 )


.param ln = 0.1u wn  = 1u

  id 0 1 100u
 xmn1 1 1 0 0 nmos1v l=ln w=wn

  vdd 2 0 1v
 xmn2 2 1 0 0 nmos1v l=ln w=wn


* vdd1  5 0 dc 5

vin1 3 0 dc 0 pulse(0 5 0ns 5ns 5ns 80ns 160ns)
vin2 4 0 dc 0 pulse(5 0 0ns 5ns 5ns 80ns 160ns)

vinA 1 0 dc 0 pulse(0 5 0ns 5ns 5ns 20ns 40ns)