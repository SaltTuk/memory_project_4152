*                1 - Input A 2 - Input B 3 - VDD 5 - Output  
.subckt nor_gate 1 2 3 5 
.param ln_nor = 0.3u wn_nor = 0.5u
.param lp_nor = 0.3u wp_nor = 1.5u

*    d g s b
xmp1 4 1 3 3 pmos1v l=lp_nor w=wp_nor
xmp2 5 2 4 3 pmos1v l=lp_nor w=wp_nor

xmn1 5 1 0 0 nmos1v l=ln_nor w=wn_nor
xmn2 5 2 0 0 nmos1v l=ln_nor w=wn_nor
.ends
