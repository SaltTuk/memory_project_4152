*                 1 - VIN 2 - VOUT  3 - VDD
.subckt not_gate 1 2 3
.param ln = 1u wn = 1u 
.param lp = 1u wp = 1u 
*    d g s b 
xmp1 2 1 3 3 pmos1v l=lp w= wp
xmn2 2 1 0 0 nmos1v l=ln w= wn

.ends