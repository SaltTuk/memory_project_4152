*                1 - Input A 2 - Input B 3 - VDD 5 - Output  
.subckt nor_gate 1 2 3 5 
.param ln = 1u wn = 1u
.param lp = 1u wp = 1u

*    d g s b
xmp1 4 1 3 3 pmos1v l=lp w= wp
xmp2 5 2 4 4 pmos1v l=lp w= wp

xmn1 5 1 0 0 nmos1v l=ln w= wn
xmn2 5 2 0 0 nmos1v l=ln w= wn
.ends
