*                R S VDD Q NQ             
.subckt sr_latch 1 2 3 4 5 
*      A B VDD OUT
xnor1  1 5 3 4 nor_gate
xnor2  2 4 3 5 nor_gate 

.ends