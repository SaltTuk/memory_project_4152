[aimspice]
[description]
234
not_gate
.include C:\Users\itsom\Desktop\FALL2022\TFE4152\90_nm_gpdk\gpdk90nm_ff.cir

.param ln = 1u wn = 1u

vdd 3 0 dc 5
vin 1 0 dc 0 pulse(0 5 10ns 1ns 1ns 25ns)
xmp1 2 1 3 3 pmos1v l=ln w= wn
xmn2 2 1 0 0 nmos1v l=ln w= wn
[dc]
1
vin
0
5
1
[tran]
0.5
50ns
X
X
0
[ana]
4 0
[end]
