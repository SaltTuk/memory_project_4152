[aimspice]
[description]
513
sr_latch
.include C:\Users\itsom\Desktop\FALL2022\TFE4152\90_nm_gpdk\gpdk90nm_ff.cir

vinA 1 0 dc 0 pulse(0 0 0ns 5ns 5ns 80ns 160ns)
vinB 2 0 dc 0 pulse(0 5 0ns 5ns 5ns 40ns 80ns)
vdd1  3 0 dc 5
vdd2  6 0 dc 5


xnor1  1 5 3 4 nor_gate
xnor2  2 4 6 5 nor_gate 

** NOR GATE     Input A , Input B , VDD, Output
.subckt nor_gate 1 2 3 5
.param ln = 1u wn = 1u

xmp1 4 1 3 3 pmos1v l=ln w= wn
xmp2 5 2 4 4 pmos1v l=ln w= wn

xmn1 5 1 0 0 nmos1v l=ln w= wn
xmn2 5 2 0 0 nmos1v l=ln w= wn
.ends

[dc]
1
vdd
0
5
0.2
[tran]
1
320ns
X
X
0
[ana]
4 5
0
1 1
1 1 -1 6
3
v(2)
v(4)
v(5)
0
1 1
1 1 -1 6
2
v(4)
v(5)
0
1 1
1 1 0 5
2
v(1)
v(2)
0
1 1
1 1 -1 6
1
v(5)
0
1 1
1 1 -1 6
1
v(4)
[end]
